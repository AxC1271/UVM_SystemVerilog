`timescale 1ns / 1ps

/*================================================
File Name: interface.sv
Description: interface description
Author: Andrew Chen
Date Created: Dec 17 2025
================================================*/

interface axi_interface();

    // input signals

    // output signals

endinterface