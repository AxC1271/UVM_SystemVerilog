`timescale 1ns / 1ps

/*================================================
File Name: axilite_slave.sv
Description: axi slave device
Author: Andrew Chen
Date Created: Dec 16 2025
================================================*/

module axilite_slave (

);

endmodule