`timescale 1ns / 1ps

/*================================================
File Name: axilite_slave.sv
Description: axi slave device (memory)
Author: Andrew Chen
Date Created: Dec 16 2025
================================================*/

module axilite_slave (
    // global
    input wire ACLK,
    input wire ARESETn
);

endmodule